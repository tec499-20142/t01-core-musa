`timescale 1ns/100ps

module modelo_referencia (xclk);

parameter XCLK_FREQ    = 48000000;

input  wire                 xclk;         


endmodule

