`timescale 1ns/100ps

module codigo (xclk);

//reg [31:0]  dados [tamanho da memoria];     

parameter   XCLK_FREQ       = 48000000;    // Frequency in Hz of xclk

input  wire                   xclk;  // external interface clock

//initial $readmemb("Estimulos.b", dados);
  

endmodule
