library verilog;
use verilog.vl_types.all;
entity modelo_tb is
end modelo_tb;
