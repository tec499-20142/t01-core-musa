library verilog;
use verilog.vl_types.all;
entity musa_monitor_sv_unit is
end musa_monitor_sv_unit;
