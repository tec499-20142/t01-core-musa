library verilog;
use verilog.vl_types.all;
entity musa_data_item_sv_unit is
end musa_data_item_sv_unit;
