library verilog;
use verilog.vl_types.all;
entity musa_tb is
end musa_tb;
