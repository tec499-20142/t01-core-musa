library verilog;
use verilog.vl_types.all;
entity opcodes_sv_unit is
end opcodes_sv_unit;
