library verilog;
use verilog.vl_types.all;
entity defines_sv_unit is
end defines_sv_unit;
