library verilog;
use verilog.vl_types.all;
entity dut_tb is
end dut_tb;
